-- File:	BRepTools_ReShape.cdl
-- Created:	Wed Jun  3 12:43:06 1998
-- Author:	data exchange team
--		<det@loufox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1998


class ReShape from BRepTools inherits TShared from MMgt

    ---Purpose: Rebuilds a Shape by making pre-defined substitutions on some
    --          of its components
    --
    --          In a first phase, it records requests to replace or remove
    --          some individual shapes
    --          For each shape, the last given request is recorded
    --          Requests may be applied "Oriented" (i.e. only to an item with
    --          the SAME orientation) or not (the orientation of replacing
    --          shape is respectful of that of the original one)
    --           
    --          Then, these requests may be applied to any shape which may
    --          contain one or more of these individual shapes
    --
    --          Requests stored in another ReShape object can be accumulated into
    --          \a this object using the Join() method.

uses 
    ShapeEnum from TopAbs, 
    Shape     from TopoDS,
    DataMapOfShapeShape from TopTools

is

    Create returns mutable ReShape from BRepTools;
    	---Purpose: Returns an empty Reshape

    Clear (me: mutable);
    	---Purpose: Clears all substitutions requests

    Remove (me: mutable; shape: Shape from TopoDS;
    	    oriented: Boolean = Standard_False);
    	---Purpose: Sets a request to Remove a Shape
    	--          If <oriented> is True, only for a shape with the SAME
    	--          orientation. Else, whatever the orientation

    Replace (me: mutable; shape, newshape: Shape from TopoDS;
    	     oriented: Boolean = Standard_False);
    	---Purpose: Sets a request to Replace a Shape by a new one
    	--          If <oriented> is True, only if the orientation is the same
    	--          Else, whatever the orientation, and the new shape takes the
    	--          same orientation as <newshape> if the replaced one has the
    	--          same as <shape>, else it is reversed

    IsRecorded (me; shape: Shape from TopoDS) returns Boolean;
	---Purpose: Tells if a shape is recorded for Replace/Remove

    Value (me; shape: Shape from TopoDS) returns Shape from TopoDS;
    	---Purpose: Returns the new value for an individual shape
    	--          If not recorded, returns the original shape itself
    	--          If to be Removed, returns a Null Shape
    	--          Else, returns the replacing item

    Status (me: mutable; shape: Shape from TopoDS; newsh: out Shape from TopoDS; last : Boolean = Standard_False)
    returns Integer is virtual;
    	---Purpose: Returns a complete substitution status for a shape
    	--          0  : not recorded,   <newsh> = original <shape>
    	--          < 0: to be removed,  <newsh> is NULL
    	--          > 0: to be replaced, <newsh> is a new item
	--          If <last> is False, returns status and new shape recorded in
	--          the map directly for the shape, if True and status > 0 then
	--          recursively searches for the last status and new shape.

    Apply (me: mutable; shape: Shape from TopoDS; until: ShapeEnum from TopAbs; buildmode: Integer)
    returns Shape from TopoDS is virtual;
    	---Purpose: Applies the substitutions requests to a shape
    	--         
    	--          <until> gives the level of type until which requests are taken
    	--          into account. For subshapes of the type <until> no rebuild 
        --          and futher exploring are done.
    	--          ACTUALLY, NOT IMPLEMENTED BELOW  TopAbs_FACE
    	--           
    	--          <buildmode> says how to do on a SOLID,SHELL ... if one of its
    	--          sub-shapes has been changed:
    	--          0: at least one Replace or Remove -> COMPOUND, else as such
    	--          1: at least one Remove (Replace are ignored) -> COMPOUND
    	--          2: Replace and Remove are both ignored
    	--          If Replace/Remove are ignored or absent, the result as same
    	--          type as the starting shape

    Apply (me: mutable; shape: Shape from TopoDS; until: ShapeEnum from TopAbs = TopAbs_SHAPE)
    returns Shape from TopoDS is virtual;
    	---Purpose: Applies the substitutions requests to a shape.
    	--         
    	--          <until> gives the level of type until which requests are taken
    	--          into account. For subshapes of the type <until> no rebuild 
        --          and futher exploring are done.
	--
	--          NOTE: each subshape can be replaced by shape of the same type
	--          or by shape containing only shapes of that type (for 
	--          example, TopoDS_Edge can be replaced by TopoDS_Edge,
	--          TopoDS_Wire or TopoDS_Compound containing TopoDS_Edges).
	--          If incompatible shape type is encountered, it is ignored
	--          and flag FAIL1 is set in Status.

    Join (me: mutable; theOther: ReShape) is virtual;
    ---Purpose: Adds mapping of \a theOther into \a this.
    --          Thus, \a this will contain a cumulative map. This can be used,
    --          for example, for concurrent shape processing and then reduction
    --          (i.e. accumulation of results in a single object).
    ---Warning: \a theOther and \a this should be consistent (e.g. they should
    --          not contain the same subshapes, or ModeConsiderLocation() and
    --          ModeConsiderOrientation() should be the same).
    
    ModeConsiderLocation(me: mutable) returns Boolean;
    ---C++: return &
    ---Purpose:Returns (modifiable) the flag which defines whether Location of shape take into account
    --         during replacing shapes.

    ModeConsiderOrientation(me: mutable) returns Boolean;
    ---C++: return &
    ---Purpose:Returns (modifiable) the flag which defines whether Orientation of shape take into account
    --         during replacing shapes.

fields

    myNMap: DataMapOfShapeShape from TopTools;  -- normal case
    myRMap: DataMapOfShapeShape from TopTools;  -- REVERSED
    myStatus: Integer is protected; -- error status
    myConsiderLocation    : Boolean;
    myConsiderOrientation : Boolean;

end ReShape;
