-- File:	ProjLib_CompProjectedCurve.cdl
-- Created:	Mon Sep 22 12:46:50 1997
-- Author:	Roman BORISOV
--		<rbv@pronox.nnov.matra-dtv.fr>
---Copyright:	 Matra Datavision 1997

class CompProjectedCurve from ProjLib inherits Curve2d  from   Adaptor2d
    
uses
    HSurface from Adaptor3d, 
    HCurve   from Adaptor3d,  
    HCurve2d   from Adaptor2d,
    Pnt2d  from  gp, 
    Vec2d  from  gp, 
    Pnt  from  gp,
    Array1OfReal   from  TColStd,  
    HSequenceOfHSequenceOfPnt  from  ProjLib,
    Shape  from  GeomAbs, 
    HArray1OfBoolean  from  TColStd, 
    HArray1OfReal  from  TColStd,
    CurveType  from  GeomAbs

raises
    
    OutOfRange          from Standard,
    NoSuchObject        from Standard,
    DomainError         from Standard,
    NotImplemented      from Standard
    
is
 
    Create  returns  CompProjectedCurve; 
     
     
    Create(S   : HSurface from Adaptor3d; 
    	   C   : HCurve   from Adaptor3d; 
    	   TolU,  TolV:  Real  from  Standard) 
    returns CompProjectedCurve; 
    ---Purpose: try to find all solutions 

    Create(S   : HSurface from Adaptor3d; 
    	   C   : HCurve   from Adaptor3d; 
    	   TolU,  TolV,  MaxDist:  Real  from  Standard) 
    returns CompProjectedCurve;  
    ---Purpose: this constructor tries to optimize the search using the 
    -- assamption that maximum distance between surface and curve less or 
    -- equal then MaxDist. 
    -- if MaxDist < 0 then algorithm works as above.
        
    Init(me:  in  out) 
    ---Purpose : computes a set of projected point and determine the 
    -- continuous parts of the projected  curves. The  points  
    -- corresponding to a projection on the bounds of the surface are  
    -- included  in this set of points.    
    is  static; 
    
    Load(me : in out;S : HSurface from Adaptor3d)
	---Purpose: Changes the surface.
    is static;
    
    Load(me : in out; C : HCurve from Adaptor3d)
	---Purpose: Changes the  curve.
    is static; 

    GetSurface(me) returns HSurface from Adaptor3d
	---C++: return const &
    is static;

    GetCurve(me) returns  HCurve from Adaptor3d 
	---C++: return const &
    is static;
   
    GetTolerance(me;  TolU,  TolV:  in  out  Real) 
    is  static;
     --
    --     Global methods - Apply to the whole curve.
    --     
    NbCurves (me) returns Integer  from  Standard
    ---Purpose: returns the number of continuous part of the projected curve
    is static;

    Bounds(me; Index : in Integer from  Standard; 
    	     Udeb,Ufin : out Real  from  Standard) 
    --- Purpose : returns the bounds of the continuous part corresponding to Index
    raises  NoSuchObject
    is static; 
    
    IsSinglePnt(me; Index:  Integer;  P :  out  Pnt2d from gp )  returns  Boolean  from  Standard 
    --- Purpose : returns  True  if  part  of  projection with  number  Index is  a  single  point  and  writes  its  coordinats in  P 
    raises  NoSuchObject
    is  static;
 
    IsUIso(me; Index:  Integer;  U :  out  Real from Standard)  returns  Boolean  from  Standard 
    --- Purpose : returns  True  if  part  of  projection with  number  Index is  an  u-isoparametric curve  of  input  surface     
    raises  NoSuchObject
    is  static;
 
    IsVIso(me; Index:  Integer;  V :  out  Real from Standard)  returns  Boolean  from  Standard 
    --- Purpose : returns  True  if  part  of  projection with  number  Index is  an  v-isoparametric curve  of  input  surface 
    raises  NoSuchObject
    is  static;


    Value(me; U : Real from  Standard) returns Pnt2d  from gp
    --- Purpose : Computes the point of parameter U on the curve.
    is  redefined  static;
    
    D0 (me; U : Real from  Standard; P : out Pnt2d from gp)
         --- Purpose : Computes the point of parameter U on the curve. 
    raises  DomainError 
    is  redefined  static;
    
    D1 (me; U : Real from  Standard; P : out Pnt2d from gp ; V : out Vec2d from gp)
         --- Purpose : Computes the point of parameter U on the curve with its
         --  first derivative.
     raises 
    	DomainError from Standard
        --- Purpose : Raised if the continuity of the current interval
        --  is not C1.

    is  redefined   static; 
     
    D2 (me; U : Real from  Standard; P : out Pnt2d from gp; V1, V2 : out Vec2d from gp)
        --- Purpose :
        --  Returns the point P of parameter U, the first and second
        --  derivatives V1 and V2.
     raises 
    	DomainError from Standard
        --- Purpose : Raised if the continuity of the current interval
        --  is not C2.
     is  redefined static; 
      
    DN (me; U : Real; N : Integer)   returns Vec2d from gp
        --- Purpose :
        --  The returned vector gives the value of the derivative for the 
        --  order of derivation N.
     raises  
        OutOfRange from Standard,
        --- Purpose : Raised if N < 1. 
        NotImplemented  from  Standard  
	--- Purpose : Raised if N > 2.

    is redefined  static; 
 
    FirstParameter(me)  returns  Real 
    	---Purpose: Returns  the  first  parameter of  the  curve  C 
	--  which  has  a  projection  on  S. 
    is  redefined  static; 
     
    LastParameter(me)  returns  Real 
    	---Purpose: Returns  the  last  parameter of  the  curve  C 
	--  which  has  a  projection  on  S. 
    is redefined  static; 

    NbIntervals(me; S : Shape from GeomAbs) returns Integer
	---Purpose: Returns  the number  of  intervals which  define   
    	--  an  S  continuous  part  of  the  projected  curve
   is  redefined  static;
 
    Trim(me;FirstParam,LastParam,Tol  :  Real)  returns HCurve2d  from  Adaptor2d
	---Purpose: Returns    a  curve equivalent   of  <me>  between
	--          parameters <First>  and <Last>. <Tol>  is used  to
	--          test for 2d points confusion.
      raises
    	OutOfRange from Standard
	---Purpose: If <First> >= <Last> 
     is redefined static;

	
    Intervals(me; T : in out Array1OfReal from TColStd; 
    	          S : Shape from GeomAbs)
	---Purpose: Returns  the  parameters  corresponding  to
	--          S  discontinuities.
	--          
	--          The array must provide  enough room to  accomodate
	--          for the parameters. i.e. T.Length() > NbIntervals()
   raises
    	OutOfRange from Standard 
   is   redefined  static;
 
    BuildIntervals(me;  S : Shape from GeomAbs)
    raises
    	OutOfRange from Standard 
    is private;
 
    MaxDistance(me;  Index:  Integer)   
        ---Purpose:  returns  the  maximum  distance  between   
    	--  curve  to  project  and  surface
    returns  Real 
    raises  NoSuchObject;
    
--  Methods  for  debugging 
    GetSequence(me) returns  HSequenceOfHSequenceOfPnt  from  ProjLib 
     ---C++: return const &
    is static; 
     
    GetType(me) returns CurveType from GeomAbs
	---Purpose: Returns  the  type of the   curve  in the  current
	--          interval :   Line,   Circle,   Ellipse, Hyperbola,
	--          Parabola, BezierCurve, BSplineCurve, OtherCurve.
    is redefined  static;
      
fields

  mySurface     :  HSurface                  from  Adaptor3d; 
  myCurve       :  HCurve                    from  Adaptor3d; 
  myNbCurves    :  Integer                   from  Standard; 
  mySequence    :  HSequenceOfHSequenceOfPnt from  ProjLib; 
  myTolU        :  Real                      from  Standard;
  myTolV        :  Real                      from  Standard; 
  myMaxDist     :  Real                      from  Standard;  
  myUIso        :  HArray1OfBoolean          from  TColStd;
  myVIso        :  HArray1OfBoolean          from  TColStd;
  mySnglPnts    :  HArray1OfBoolean          from  TColStd;    
  myMaxDistance :  HArray1OfReal             from  TColStd; 
  TabInt        :  HArray1OfReal             from  TColStd;
        
end CompProjectedCurve;
