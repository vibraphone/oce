-- File:	Approx_ComputeLine.cdl
-- Created:	Tue Jan 26 11:50:18 1993
-- Author:	Laurent PAINNOT
--		<lpa@sdsun1>
---Copyright:	 Matra Datavision 1993



generic class ComputeLine from Approx 
    	    	    (MultiLine as any;
    	    	     LineTool  as any) --as TheLineTool(MultiLine)


uses ParametrizationType       from Approx,
     SequenceOfReal            from TColStd,
     HArray1OfReal             from TColStd,
     Array1OfReal              from TColStd,
     SequenceOfMultiCurve      from AppParCurves,
     HArray1OfMultiCurve       from AppParCurves,
     HArray1OfConstraintCouple from AppParCurves,
     Constraint                from AppParCurves,
     SequenceOfHArray1OfReal   from Approx,
     MultiCurve                from AppParCurves,
     MultiBSpCurve             from AppParCurves,
     Vector                    from math
     
     

private class MyGradient instantiates Gradient from AppParCurves
    	    	    	    	       (MultiLine,
			    	    	LineTool);
							  
is


    Create(Line:            MultiLine; 
    	   degreemin:       Integer = 4;
           degreemax:       Integer = 8;
    	   Tolerance3d:     Real    = 1.0e-3; 
    	   Tolerance2d:     Real    = 1.0e-6;
           NbIterations:    Integer = 5;
	   cutting:         Boolean = Standard_True; 
    	   parametrization: ParametrizationType from Approx =
    	   Approx_ChordLength;
	   Squares:         Boolean = Standard_False)
	   
	---Purpose: The MultiLine <Line> will be approximated until tolerances
	--          will be reached.
	--          The approximation will be done from degreemin to degreemax
	--          with a cutting if the corresponding boolean is True.
	--          If <Squares> is True, the computation will be done with
	--          no iteration at all.

    returns ComputeLine;


    Create(Line:         MultiLine; 
    	   Parameters:   Vector from math;
    	   degreemin:    Integer = 4;
    	   degreemax:    Integer = 8;
    	   Tolerance3d:  Real    = 1.0e-03; 
    	   Tolerance2d:  Real    = 1.0e-06; 
	   NbIterations: Integer = 5;
	   cutting:      Boolean = Standard_True; 
    	   Squares:      Boolean = Standard_False)
	   
	---Purpose: The MultiLine <Line> will be approximated until tolerances
	--          will be reached.
	--          The approximation will be done from degreemin to degreemax
	--          with a cutting if the corresponding boolean is True.
	--          If <Squares> is True, the computation will be done with
	--          no iteration at all.

    returns ComputeLine;


    Create(Parameters:   Vector from math;
    	   degreemin:    Integer = 4;
    	   degreemax:    Integer = 8;
    	   Tolerance3d:  Real    = 1.0e-03; 
    	   Tolerance2d:  Real    = 1.0e-06; 
	   NbIterations: Integer = 5;
	   cutting:      Boolean = Standard_True; 
    	   Squares:      Boolean = Standard_False)
	   
	---Purpose: Initializes the fields of the algorithm.

    returns ComputeLine;


    Create(degreemin:    Integer = 4;
    	   degreemax:    Integer = 8;
    	   Tolerance3d:  Real    = 1.0e-03; 
    	   Tolerance2d:  Real    = 1.0e-06; 
	   NbIterations: Integer = 5;
	   cutting:      Boolean = Standard_True; 
    	   parametrization: ParametrizationType from Approx =
    	   Approx_ChordLength;
    	   Squares:      Boolean = Standard_False)
	   
	---Purpose: Initializes the fields of the algorithm.

    returns ComputeLine;


    Init(me: in out; degreemin:    Integer = 4;
    	             degreemax:    Integer = 8;
    	             Tolerance3d:  Real    = 1.0e-03; 
    	             Tolerance2d:  Real    = 1.0e-06; 
	             NbIterations: Integer = 5;
	             cutting:      Boolean = Standard_True; 
    	             parametrization: ParametrizationType from Approx =
    	             Approx_ChordLength;
    	             Squares:      Boolean = Standard_False)
	   
	---Purpose: Initializes the fields of the algorithm.

    is static;




    Perform(me: in out; Line: MultiLine)
	---Purpose: runs the algorithm after having initialized the fields.
    
    is static;


    Compute(me: in out; Line: MultiLine; fpt, lpt: Integer;
    	    Para: in out Vector from math; TheTol3d, TheTol2d: in out Real)
	---Purpose: is internally used in the algorithm.

    returns Boolean
    is static private;
    
    
    ComputeCurve(me: in out; Line: MultiLine; firspt, lastpt: Integer) 
	---Purpose: is internally used in the algorithm.
    
    returns Boolean
    is static private;
    
    
    Parameters(me; Line: MultiLine; firstP, LastP: Integer;
               TheParameters: in out Vector)
    	---Purpose: computes new parameters between firstP and lastP.

    is static private;
    
    
    SetDegrees(me: in out; degreemin, degreemax: Integer)
    	---Purpose: changes the degrees of the approximation.
    
    is static;
    
    
    SetTolerances(me: in out; Tolerance3d, Tolerance2d: Real)
    	---Purpose: Changes the tolerances of the approximation.
    
    is static;
    

    SetConstraints(me: in out; firstC, lastC: Constraint from AppParCurves)
    	    ---Purpose: changes the first and the last constraint points.
    is static;


    IsAllApproximated(me) 
    	---Purpose: returns False if at a moment of the approximation,
    	--          the status NoApproximation has been sent by the user
    	--          when more points were needed.
    
    returns Boolean
    is static;
    

    IsToleranceReached(me)
    	---Purpose: returns False if the status NoPointsAdded has been sent.
    
    returns Boolean
    is static;
    

    Error(me; Index: Integer; tol3d: in out Real; tol2d: in out Real)
    	---Purpose: returns the tolerances 2d and 3d of the <Index> MultiCurve.

    is static;
    

    NbMultiCurves(me)
    	---Purpose: Returns the number of MultiCurve doing the approximation
    	--          of the MultiLine.
    returns Integer
    is static;


    Value(me; Index: Integer = 1)
    	---Purpose: returns the result of the approximation.
    	---C++: return const&
    returns MultiCurve from AppParCurves
    is static;

    ChangeValue(me: in out; Index: Integer = 1)
    	---Purpose: returns the result of the approximation.
    	---C++: return &
    returns MultiCurve from AppParCurves
    is static;


    SplineValue(me: in out)
    	---Purpose: returns the result of the approximation.
    	---C++: return const&
    returns MultiBSpCurve from AppParCurves
    is static;

    Parametrization(me; partype :  in  out ParametrizationType from Approx) 
    	---Purpose: returns the type  of  parametrization
    is static;


    Parameters(me; Index: Integer = 1)
    	---Purpose: returns the new parameters of the approximation
    	--          corresponding to the points of the multicurve <Index>.
    	---C++: return const&
    returns Array1OfReal from TColStd
    is static;
 
     
    
    SearchFirstLambda(me; Line: MultiLine; Para: Vector; 
    	    	      V: Vector; index: Integer)
    returns Real
    is static private;
    
    SearchLastLambda(me: ; Line: MultiLine; Para: Vector;
    	    	     V: Vector; index: Integer)
    returns Real
    is static private;
    
    FirstTangencyVector(me; Line: MultiLine; index: Integer; V: in out Vector)
    is static private;
    
    LastTangencyVector(me; Line: MultiLine; index: Integer; V: in out Vector)
    is static private;


fields


myMultiCurves: SequenceOfMultiCurve      from AppParCurves;    
TheMultiCurve: MultiCurve                from AppParCurves;
myspline     : MultiBSpCurve             from AppParCurves;
alldone:       Boolean                   from Standard;
tolreached:    Boolean                   from Standard;
Par:           ParametrizationType       from Approx;
myParameters:  HArray1OfReal             from TColStd;
myfirstParam:  HArray1OfReal             from TColStd;
myPar:         SequenceOfHArray1OfReal   from Approx;
Tolers3d:      SequenceOfReal            from TColStd;
Tolers2d:      SequenceOfReal            from TColStd;
myConstraints: HArray1OfConstraintCouple from AppParCurves;
mydegremin:    Integer                   from Standard;
mydegremax:    Integer                   from Standard;
mytol3d:       Real                      from Standard;
mytol2d:       Real                      from Standard;
currenttol3d:  Real                      from Standard;
currenttol2d:  Real                      from Standard;
mycut:         Boolean                   from Standard;
mysquares:     Boolean                   from Standard;
myitermax:     Integer                   from Standard;
myfirstC:      Constraint                from AppParCurves;
mylastC:       Constraint                from AppParCurves;
IsClear:       Boolean                   from Standard;
nbML:          Integer                   from Standard;

end ComputeLine;
